/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_mixcol.v                                                               *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Testbench block AES - 128 bit input, s-box 4 BRAM, 3 cycle round                              *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

`timescale 1ns / 1ps

module aes_128_mixcol_tb;

 /*************************************************************************************
 *            PARAMETERS                                                             *
 *************************************************************************************/
parameter clk_dly = 20;

/*************************************************************************************
 *            INTERNAL WIRES & REGS                                                  *
 *************************************************************************************/
//inputs
reg		clk;
reg		en;
reg	[127:0]	in_data;

//output
wire	[127:0]	out_data;

 /*************************************************************************************
 *            BLOCK INSTANCE                                                          *
 *************************************************************************************/
aes_128_mixcol aes_128_mixcol (		.clk(clk),
					.en(en),
					.in_data(in_data),
					.out_data(out_data));

/*************************************************************************************
 *            INITIAL                                                                *
 *************************************************************************************/
//initialization clock signals
initial
begin
	clk = 1'b0;
end

always
#clk_dly clk = ~clk;

//initial full
initial
begin
	wait_n_clocks(3);
	aes_128_mixcol_ini;
	aes_128_mixcol_set_data;
end

/*************************************************************************************
 *            TASKS                                                                  *
 *************************************************************************************/
//initialization all signal
task aes_128_mixcol_ini;
begin
	en = 1'b0;
	in_data = 128'b0;
end
endtask

/**************************************************************************************************/
// wait N clocks

task wait_n_clocks;
input integer N;
integer n; 
begin
	@(posedge clk);
	for (n = 0; n < N; n = n + 1)
		@(posedge clk);
end
endtask

/**************************************************************************************************/
//set data
task aes_128_mixcol_set_data;
begin
	@(posedge clk);
	//in_data <= 128'h876e46a6f24ce78c4d904ad897ecc395;
	in_data <= 128'he7d0caba51b770cd04e160098ce05363;
	@(posedge clk);
	en <= 1'b1;
	in_data <= 128'he7d0caba51b770cd04e160098ce05363;
	@(posedge clk);
	en <= 1'b0;
	in_data <= 128'b0;
end
endtask

/**************************************************************************************************/

endmodule
