/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_core.v                                                                 *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Block AES - 128 bit input, s-box 4 BRAM, 3 cycle round                                        *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

module aes_128_core (
	clk,
	kill,
	en_mixcol,
	start,
	rounds_end,
	in_data,
	key_round,

	out_data
	);

/**************************************************************************************************
*        I/O PORTS
 **************************************************************************************************/
input			clk;
input			kill;
input			en_mixcol;
input			start;
input			rounds_end;
input	[127:0]		in_data;
input	[127:0]		key_round;

output	[127:0]		out_data;

/**************************************************************************************************
 *      LOCAL WIRES, REGS                                                                         *
 **************************************************************************************************/
wire	[127:0]		mixcol_out;
wire	[127:0]		subbytes_out;

reg	[127:0]		round_data;

/**************************************************************************************************
 *      LOGIC                                                                                     *
 **************************************************************************************************/
//SubBytes and ShiftRows
aes_128_subbytes aes_128_subbytes (	.clk(clk),
					.kill(kill),
					.en(1'b1),
					.in_data(round_data),
					.out_data(subbytes_out));

/**************************************************************************************************/
//MixColums
aes_128_mixcol aes_128_mixcol (		.clk(clk),
					.kill(kill),
					.en(en_mixcol),
					.in_data(subbytes_out),
					.out_data(mixcol_out));

/**************************************************************************************************/
//AddRoundKey
always @(posedge clk)
	if (kill)
		round_data <= 128'b0;
	else if (start)
		round_data <= in_data ^ key_round;
	else
		round_data <= mixcol_out ^ key_round;

/**************************************************************************************************/
//Output data
assign out_data = (rounds_end) ? round_data : 128'b0;

/**************************************************************************************************/

endmodule







