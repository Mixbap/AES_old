/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_subbytes_tb.v                                                          *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Block AES - 128 bit input, s-box 4 BRAM, 3 cycle round                                        *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

`timescale 1ns / 1ps

module aes_128_subbytes_tb;

 /*************************************************************************************
 *            PARAMETERS                                                             *
 *************************************************************************************/
parameter clk_dly = 20;
parameter rst_dly = 50;

/*************************************************************************************
 *            INTERNAL WIRES & REGS                                                  *
 *************************************************************************************/
//inputs
reg		clk;
reg		kill;
reg		en;
reg	[127:0]	in_data;

//output
wire	[127:0]	out_data;

 /*************************************************************************************
 *            BLOCK INSTANCE                                                          *
 *************************************************************************************/
aes_128_subbytes aes_128_subbytes (	.clk(clk),
					.kill(kill),
					.en(en),
					.in_data(in_data),
					.out_data(out_data));

/*************************************************************************************
 *            INITIAL                                                                *
 *************************************************************************************/
//initialization clock signals
initial
begin
	clk = 1'b0;
	kill = 1'b0;
end

always
#clk_dly clk = ~clk;

//initial full
initial
begin
	aes_128_subbytes_rst;
	aes_128_subbytes_ini;
	wait_n_clocks(3);
	aes_128_subbytes_set_data;
end

/*************************************************************************************
 *            TASKS                                                                  *
 *************************************************************************************/
//reset signal
task aes_128_subbytes_rst;
begin
	kill <= 1'b1;
	#rst_dly kill <= 1'b0;
end
endtask

/**************************************************************************************************/
//initialization all signal
task aes_128_subbytes_ini;
begin
	en = 0;
	in_data = 128'b0;
end
endtask

/**************************************************************************************************/
// wait N clocks

task wait_n_clocks;
input integer N;
integer n; 
begin
	@(posedge clk);
	for (n = 0; n < N; n = n + 1)
		@(posedge clk);
end
endtask

/**************************************************************************************************/
//set data
task aes_128_subbytes_set_data;
begin
	@(posedge clk);
	en <= 1'b1;
	in_data <= 128'hf0e0d0c0b0a090807060504030201000;
	@(posedge clk);
	en <= 1'b0;
	in_data <= 128'b0;
end
endtask
/**************************************************************************************************/

endmodule
