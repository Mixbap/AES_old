/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_keyram_2key.v                                                          *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Block AES - 128 bit input, s-box 4 BRAM, 4 cycle round                                        *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

(* keep_hierarchy = "yes" *)

module aes_128_keyram_2key (
	/* inputs */
	input			clk,
	input			kill,
	input			en_wr,
	input		[63:0]	key_round_wr,
	input			key_ready,
	
	/* outputs */
	output		[127:0]	key_round_rd,
	output			wr_idle
	);

/**************************************************************************************************
 *      LOCAL WIRES, REGS                                                                         *
 **************************************************************************************************/
wire		[63:0]	ram_out;
wire		[5:0]	addr_wr;
wire		[5:0]	addr_rd;

/**************************************************************************************************
 *      LOGIC                                                                                     *
 **************************************************************************************************/
aes_128_keyram_mem_2key aes_128_keyram_mem_2key(	.clk(clk),
							.kill(kill),
							.en_wr(en_wr),
							.addr_wr(addr_wr),
							.addr_rd(addr_rd),
							.key_round_wr(key_round_wr),
							.ram_out(ram_out));

/**************************************************************************************************/					
aes_128_keyram_control_2key aes_128_keyram_control_2key(.clk(clk),
							.kill(kill),
							.en_wr(en_wr),
							.key_ready(key_ready),
							.ram_out(ram_out),
							.key_round_rd(key_round_rd),
							.addr_wr(addr_wr),
							.addr_rd(addr_rd),
							.wr_idle(wr_idle));

/**************************************************************************************************/
endmodule







