/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_sbox_tb.v                                                              *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Testbench block AES - 128 bit input, s-box 4 BRAM, 3 cycle round                              *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

`timescale 1ns / 1ps

module aes_128_sbox_tb;

 /*************************************************************************************
 *            PARAMETERS                                                             *
 *************************************************************************************/
parameter clk_dly = 20;

/*************************************************************************************
 *            INTERNAL WIRES & REGS                                                  *
 *************************************************************************************/
//inputs
reg		clk;
reg	[7:0]	addra;
reg	[7:0]	addrb;

//outputs
wire	[7:0]	doa;
wire	[7:0]	dob;

 /*************************************************************************************
 *            BLOCK INSTANCE                                                          *
 *************************************************************************************/
aes_128_sbox aes_128_sbox(		.clka(clk),
					.clkb(clk),
					.wea(1'b0),
					.web(1'b0),
					.addra(addra),
					.addrb(addrb),
					.dia(),
					.dib(),
					.doa(doa),
					.dob(dob));

/*************************************************************************************
 *            INITIAL                                                                *
 *************************************************************************************/
//initialization clock signals
initial
begin
	clk = 1'b0;
end

always
#clk_dly clk = ~clk;

//initial full
initial
begin
	wait_n_clocks(3);
	aes_128_sbox_ini;
	aes_128_sbox_addr;
end

/*************************************************************************************
 *            TASKS                                                                  *
 *************************************************************************************/
//initialization all signal
task aes_128_sbox_ini;
begin
	addra = 8'b0;
	addrb = 8'b0;
end
endtask

/**************************************************************************************************/
// wait N clocks

task wait_n_clocks;
input integer N;
integer n; 
begin
	@(posedge clk);
	for (n = 0; n < N; n = n + 1)
		@(posedge clk);
end
endtask

/**************************************************************************************************/
//addr
task aes_128_sbox_addr;
integer i;
begin
	@(posedge clk);
	for (i = 0; i < 256; i = i + 1)
	begin
		addra <= addra + 1;
		addrb <= addrb + 1;
		@(posedge clk);
	end
end
endtask

/**************************************************************************************************/

endmodule
