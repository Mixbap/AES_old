/**************************************************************************************************
 *                                                                                                *
 *  File Name:     aes_128_key_ram.v                                                              *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:                                                                                  *
 *                                                                                                *
 *  Block AES - 128 bit input, s-box 4 BRAM, 3 cycle round                                        *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog code                                                                                  *
 **************************************************************************************************/

(* keep_hierarchy = "yes" *)

module aes_128_keyram (
	/* inputs */
	input			clk,
	input			kill,
	input			en_wr,
	input		[63:0]	key_round_wr,
	input		[4:0]	addr_wr,
	input			key_ready,
	
	/* outputs */
	output		[127:0]	key_round_rd
	);

/**************************************************************************************************
 *      LOCAL WIRES, REGS                                                                         *
 **************************************************************************************************/
wire		[63:0]	ram_out;
wire		[4:0]	addr;

/**************************************************************************************************
 *      LOGIC                                                                                     *
 **************************************************************************************************/
aes_128_keyram_mem aes_128_keyram_mem(		.clk(clk),
						.kill(kill),
						.en_wr(en_wr),
						.addr(addr),
						.key_round_wr(key_round_wr),
						.ram_out(ram_out));

/**************************************************************************************************/					
aes_128_keyram_control aes_128_keyram_control(	.clk(clk),
						.kill(kill),
						.en_wr(en_wr),
						.addr_wr(addr_wr),
						.key_ready(key_ready),
						.ram_out(ram_out),
						.key_round_rd(key_round_rd),
						.addr(addr));

/**************************************************************************************************/
endmodule







